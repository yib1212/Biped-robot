module light(
output [7:0]LED);

assign LED[7:0] = 8'b11111111;
endmodule

